`default_nettype none
module ftoi (
    input wire [31:0] x,
    output wire [31:0] y,
    input wire clk,
    input wire rstn);

wire s = x[31];
wire [7:0] e = x[30:23];
wire [22:0] m = x[22:0];
wire [31:0] absy;
//wire [23:0] rman = {1'b1, m};

assign absy =  (e < 8'b01111111) ? 32'b0 :
            (e == 8'b01111111) ? 32'b1 :
            (e == 8'b10000000) ? {31'b1, m[22]} :
            (e == 8'b10000001) ? {30'b1, m[22:21]} :
            (e == 8'b10000010) ? {29'b1, m[22:20]} :
            (e == 8'b10000011) ? {28'b1, m[22:19]} :
            (e == 8'b10000100) ? {27'b1, m[22:18]} :
            (e == 8'b10000101) ? {26'b1, m[22:17]} :
            (e == 8'b10000110) ? {25'b1, m[22:16]} :
            (e == 8'b10000111) ? {24'b1, m[22:15]} :
            (e == 8'b10001000) ? {23'b1, m[22:14]} :
            (e == 8'b10001001) ? {22'b1, m[22:13]} :
            (e == 8'b10001010) ? {21'b1, m[22:12]} :
            (e == 8'b10001011) ? {20'b1, m[22:11]} :
            (e == 8'b10001100) ? {19'b1, m[22:10]} :
            (e == 8'b10001101) ? {18'b1, m[22:9]} :
            (e == 8'b10001110) ? {17'b1, m[22:8]} :
            (e == 8'b10001111) ? {16'b1, m[22:7]} :
            (e == 8'b10010000) ? {15'b1, m[22:6]} :
            (e == 8'b10010001) ? {14'b1, m[22:5]} :
            (e == 8'b10010010) ? {13'b1, m[22:4]} :
            (e == 8'b10010011) ? {12'b1, m[22:3]} :
            (e == 8'b10010100) ? {11'b1, m[22:2]} :
            (e == 8'b10010101) ? {10'b1, m[22:1]} :
            (e == 8'b10010110) ? {9'b1, m[22:0]} :
            (e == 8'b10010111) ? {8'b1, m[22:0], 1'b0} :
            (e == 8'b10011000) ? {7'b1, m[22:0], 2'b0} :
            (e == 8'b10011001) ? {6'b1, m[22:0], 3'b0} :
            (e == 8'b10011010) ? {5'b1, m[22:0], 4'b0} :
            (e == 8'b10011011) ? {4'b1, m[22:0], 5'b0} :
            (e == 8'b10011100) ? {3'b1, m[22:0], 6'b0} :
            (e == 8'b10011101) ? {2'b1, m[22:0], 7'b0} :
            (e == 8'b10011110) ? {1'b1, m[22:0], 8'b0} : {1'b1, 31'b0};

assign y = (s == 0) ? absy : (~absy) + 1'b1;

endmodule
`default_nettype wire