`default_nettype none
module ftoi (
    input wire [31:0] x,
    output wire [31:0] y,
    input wire clk,
    input wire rstn);

wire s = x[31];     // 答えのsignビットはxの正負=x[31]に一致。
//wire [7:0] e;
//wire [22:0] m;
wire [31:0] absx = (s == 0) ? x : (~x) + 1'b1;      // 負の最大値1000...0の時に1000...0になることに注意。

assign y =  (absx[30] == 1) ? {s, 8'b10011101, absx[29:7]} + absx[6] :
            (absx[29] == 1) ? {s, 8'b10011100, absx[28:6]} + absx[5] :
            (absx[28] == 1) ? {s, 8'b10011011, absx[27:5]} + absx[4] :
            (absx[27] == 1) ? {s, 8'b10011010, absx[26:4]} + absx[3] :
            (absx[26] == 1) ? {s, 8'b10011001, absx[25:3]} + absx[2] :
            (absx[25] == 1) ? {s, 8'b10011000, absx[24:2]} + absx[1] :
            (absx[24] == 1) ? {s, 8'b10010111, absx[23:1]} + absx[0] :
            (absx[23] == 1) ? {s, 8'b10010110, absx[22:0]} :
            (absx[22] == 1) ? {s, 8'b10010101, absx[21:0], 1'b0} :
            (absx[21] == 1) ? {s, 8'b10010100, absx[20:0], 2'b0} :
            (absx[20] == 1) ? {s, 8'b10010011, absx[19:0], 3'b0} :
            (absx[19] == 1) ? {s, 8'b10010010, absx[18:0], 4'b0} :
            (absx[18] == 1) ? {s, 8'b10010001, absx[17:0], 5'b0} :
            (absx[17] == 1) ? {s, 8'b10010000, absx[16:0], 6'b0} :
            (absx[16] == 1) ? {s, 8'b10001111, absx[15:0], 7'b0} :
            (absx[15] == 1) ? {s, 8'b10001110, absx[14:0], 8'b0} :
            (absx[14] == 1) ? {s, 8'b10001101, absx[13:0], 9'b0} :
            (absx[13] == 1) ? {s, 8'b10001100, absx[12:0], 10'b0} :
            (absx[12] == 1) ? {s, 8'b10001011, absx[11:0], 11'b0} :
            (absx[11] == 1) ? {s, 8'b10001010, absx[10:0], 12'b0} :
            (absx[10] == 1) ? {s, 8'b10001001, absx[9:0], 13'b0} :
            (absx[9] == 1) ? {s, 8'b10001000, absx[8:0], 14'b0} :
            (absx[8] == 1) ? {s, 8'b10000111, absx[7:0], 15'b0} :
            (absx[7] == 1) ? {s, 8'b10000110, absx[6:0], 16'b0} :
            (absx[6] == 1) ? {s, 8'b10000101, absx[5:0], 17'b0} :
            (absx[5] == 1) ? {s, 8'b10000100, absx[4:0], 18'b0} :
            (absx[4] == 1) ? {s, 8'b10000011, absx[3:0], 19'b0} :
            (absx[3] == 1) ? {s, 8'b10000010, absx[2:0], 20'b0} :
            (absx[2] == 1) ? {s, 8'b10000001, absx[1:0], 21'b0} :
            (absx[1] == 1) ? {s, 8'b10000000, absx[0], 22'b0} :
            (absx[0] == 1) ? {s, 8'b01111111, 23'b0} : 
            (absx[31] == 1) ? {1'b1, 8'b10011110, 23'b0} : 32'b0;

endmodule
`default_nettype wire